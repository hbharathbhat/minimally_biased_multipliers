module approx_multi (a, b, r);
parameter K = 6;
parameter N = 16;
parameter M = 16;
input [N-1:0] a;
input [M-1:0] b;
output [(N+M)-1:0] r;
wire [K-3:0] m;
wire [K-3:0] n;
wire [N-1:0] l1;
wire [M-1:0] l2;
wire [(K*2)-1:0] tmp;
wire [$clog2(N)-1:0] k1;
wire [$clog2(M)-1:0] k2;
wire [$clog2(M)-1:0] p;
wire [$clog2(M)-1:0] q;
wire [$clog2(M):0] sum;
wire [K-1:0] mm;
wire [K-1:0] nn;
detect_1 #(K, N) u1(.input_a(a),.output_a(l1));
detect_1 #(K, M) u2(.input_a(b),.output_a(l2));
priorityencoder #(K, N) u3(.input_a(l1), .output_a(k1));
priorityencoder #(K, M) u4(.input_a(l2), .output_a(k2));
multiplexer #(K, N) u5(.input_a(a), .sel_line(k1), .out(m));
multiplexer #(K, M) u6(.input_a(b), .sel_line(k2), .out(n));
assign p=(k1>(K-1))?k1-(K-1):0;
assign q=(k2>(K-1))?k2-(K-1):0;
assign mm=(k1>K-1)?({1'b1,m,1'b1}):a[K-1:0];
assign nn=(k2>K-1)?({1'b1,n,1'b1}):b[K-1:0];
assign tmp=nn*mm;
assign sum=q+p;
barrelshifter #(K, N, M) u7(.input_a(tmp), .count(sum), .output_a(r));
endmodule